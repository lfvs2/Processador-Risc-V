`timescale 1ns / 1ps

module datamemory #(
    parameter DM_ADDRESS = 9,
    parameter DATA_W = 32
) (
    input logic clk,
    input logic MemRead,  // comes from control unit
    input logic MemWrite,  // comes from control unit
    input logic [DM_ADDRESS - 1:0] a,  // Read / Write address - 9 LSB bits of the ALU output
    input logic [DATA_W - 1:0] wd,  // Write Data
    input logic [2:0] Funct3,  // bits 12 to 14 of the instruction
    output logic [DATA_W - 1:0] rd  // Read Data
);

  logic [31:0] raddress;
  logic [31:0] waddress;
  logic [31:0] Datain;
  logic [31:0] Dataout;
  logic [ 3:0] Wr;

  Memoria32Data mem32 (
      .raddress(raddress),
      .waddress(waddress),
      .Clk(~clk),
      .Datain(Datain),
      .Dataout(Dataout),
      .Wr(Wr)
  );

  always_ff @(*) begin
    raddress = {{22{1'b0}}, a};
    waddress = {{22{1'b0}}, {a[8:2], {2{1'b0}}}};
    Datain = wd;
    Wr = 4'b0000;

    if (MemRead) begin // reading data functions
      case (Funct3)
        3'b000:	 // LB
            rd = {{24{Dataout[7]}}, Dataout[7:0]}; // function reads the byte with sign extension
        3'b001:  // LH
            rd = {{16{Dataout[15]}}, Dataout[15:0]} // reads half-word (16 bits) with sign extension
        3'b010:  // LW
            rd = Dataout; // reads the entire word
        3'b100:  // LBU
            rd = {24'b0, Dataout[7:0]}; // reads byte unsigned
        default: rd = Dataout; // in case of funct3 values unrecognizeds, returns the full word 
      endcase
    end else if (MemWrite) begin
      case (Funct3)
        3'b000: // SB (Store Byte)
            Wr = 4'b0001; // write byte
        3'b001: // SH (Store Half-word)
            Wr = 4'b0011; // write half-word
        3'b010: begin // SW (Store Word)
          Wr <= 4'b1111; 
          Datain <= wd;  
          end
          default: begin
          Wr <= 4'b1111;
          Datain <= wd; 
          end
         endcase
        end
    end

endmodule
